`define OP_ADD 4'b0001 // Add
`define OP_SUB 4'b0010 // Subtract
`define OP_SHL 4'b0101 // Shift Left
`define OP_SHAR 4'b0110 // Arithmetic Shift Right 
`define OP_SHLR 4'b0111 // Logical Shift Right
`define OP_RL 4'b1000 // Rotate Left
`define OP_RR 4'b1001 // Rotate Right
`define OP_AND 4'b1011 // AND
`define OP_OR 4'b1100 // OR
`define OP_XOR 4'b1101 // XOR
`define OP_NOT 4'b1110 // NOT
`define OP_MUL 4'b1111 // Multiply


module test_ALU;
	